`timescale 1ns / 1ps
//////////////////////////////////////////////////////////////////////////////////
// Company: 
// Engineer: 
// 
// Create Date: 11/06/2017 01:19:57 PM
// Design Name: 
// Module Name: high_pass_filter
// Project Name: 
// Target Devices: 
// Tool Versions: 
// Description: 
// 
// Dependencies: 
// 
// Revision:
// Revision 0.01 - File Created
// Additional Comments:
// 
//////////////////////////////////////////////////////////////////////////////////


module high_pass_filter(
    input clock,
    input ready,
    input reset,
    input coeff,
    input enable,
    input audio_in,
    output audio_out
    );
endmodule
