`timescale 1ns / 1ps
//////////////////////////////////////////////////////////////////////////////////
// Company: 
// Engineer: 
// 
// Create Date: 11/06/2017 01:19:57 PM
// Design Name: 
// Module Name: low_pass_filter
// Project Name: 
// Target Devices: 
// Tool Versions: 
// Description: 
// 
// Dependencies: 
// 
// Revision:
// Revision 0.01 - File Created
// Additional Comments:
// 
//////////////////////////////////////////////////////////////////////////////////


module low_pass_filter(
    input clock,
    input enable,
    input audio_in,
    input ready,
    output audio_out,
    input reset,
    input coeffs
    );
endmodule
